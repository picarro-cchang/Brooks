----------------------------------------------------------------------------------
-- Company:        Picarro, Inc
-- Engineer:       Sze Tan
--
-- Create Date:    04/29/2009
-- Design Name:
-- Module Name:    top_block - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all;
use work.pck_myhdl_06.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity top_block is
    port (
           clk              : in std_logic;

           rd_adc           : in unsigned(15 downto 0);
           rd_adc_clk       : out std_logic;
           rd_adc_oe        : out std_logic;

           dsp_emif_we      : in std_logic;
           dsp_emif_re      : in std_logic;
           dsp_emif_oe      : in std_logic;
           dsp_emif_ardy    : out std_logic;

           dsp_emif_ea      : in unsigned(19 downto 0);
           dsp_emif_din     : in unsigned(31 downto 0);
           dsp_emif_dout    : out unsigned(31 downto 0);

           usb_connected    : in std_logic;
           cyp_reset        : out std_logic;
           cyp_pc           : in unsigned(7 downto 0);
           dsp_ext_int4     : out std_logic;
           dsp_ext_int5     : out std_logic;
           dsp_ext_int6     : out std_logic;
           dsp_ext_int7     : out std_logic;

           dsp_clkout2      : in std_logic;
           dsp_clkout3      : in std_logic;
           dsp_eclkout      : in std_logic;

           dsp_emif_be      : in unsigned(3 downto 0);
           dsp_emif_ce      : in unsigned(3 downto 0);

           dsp_tinp0        : out std_logic;
           dsp_tinp1        : out std_logic;
           dsp_tout0        : in std_logic;
           dsp_tout1        : in std_logic;

           fp_lcd           : out unsigned(7 downto 0);
           fp_pb            : in std_logic;
           fp_rs_n          : in std_logic;
           fp_led           : out unsigned(3 downto 0);

           pwr_din          : out unsigned(7 downto 0);
           pwr_dout         : in unsigned(7 downto 0);

           aux_din          : out unsigned(3 downto 0);
           aux_dout         : in unsigned(3 downto 0);

           monitor          : out std_logic;

           lsr1_sck         : out std_logic;
           lsr1_ss          : out std_logic;
           lsr1_rd          : out std_logic;
           lsr1_mosi        : out std_logic;
           lsr1_disable     : out std_logic;

           lsr2_sck         : out std_logic;
           lsr2_ss          : out std_logic;
           lsr2_rd          : out std_logic;
           lsr2_mosi        : out std_logic;
           lsr2_disable     : out std_logic;

           lsr3_sck         : out std_logic;
           lsr3_ss          : out std_logic;
           lsr3_rd          : out std_logic;
           lsr3_mosi        : out std_logic;
           lsr3_disable     : out std_logic;

           lsr4_sck         : out std_logic;
           lsr4_ss          : out std_logic;
           lsr4_rd          : out std_logic;
           lsr4_mosi        : out std_logic;
           lsr4_disable     : out std_logic;

           wmm_refl1        : in std_logic;
           wmm_refl2        : in std_logic;
           wmm_tran1        : in std_logic;
           wmm_tran2        : in std_logic;
           wmm_busy1        : in std_logic;
           wmm_busy2        : in std_logic;
           wmm_rd           : out std_logic;
           wmm_convst       : out std_logic;
           wmm_clk          : out std_logic;

           sw1              : out std_logic;
           sw2              : out std_logic;
           sw3              : out std_logic;
           sw4              : out std_logic;

           lsr1_0           : out std_logic;
           lsr1_1           : out std_logic;
           lsr2_0           : out std_logic;
           lsr2_1           : out std_logic;
           lsr3_0           : out std_logic;
           lsr3_1           : out std_logic;
           lsr4_0           : out std_logic;
           lsr4_1           : out std_logic;

           mictor           : out unsigned(33 downto 0);
           fpga_led         : out unsigned(3 downto 0);

           i2c_rst0         : out std_logic;
           i2c_rst1         : out std_logic;

           i2c_scl0         : in std_logic;
           i2c_sda0         : in std_logic;
           i2c_scl1         : in std_logic;
           i2c_sda1         : in std_logic
    );
end top_block;

architecture behavioral of top_block is
begin
    dsp_emif_ardy <= '0';
end behavioral;
